`timescale 1ns / 1ps

// =============================================================
// dm: 数据存储器 (Data Memory) - 256 字节 RAM
// =============================================================
// 功能: 实现 CPU 的数据存储器，支持多种访存宽度
//
// 设计要点:
// - mem[] 是 8 位宽 (1 字节) 的数组，按"字节寻址"
// - addr 每 +1 表示下一个字节
// - 读数据: 组合逻辑 always @(*)，根据 DMType 拼出 32 位 dout
// - 写数据: 时序逻辑 always @(posedge clk)，DMWr=1 时写入
// =============================================================

// =============================================================
// DMType/Funct3 编码对照表
// =============================================================
// DMType | Load指令 | Store指令 | 访问宽度 | 扩展方式
// -------|----------|-----------|----------|----------
// 3'b000 | LB       | SB        | 8-bit    | 符号扩展
// 3'b001 | LH       | SH        | 16-bit   | 符号扩展
// 3'b010 | LW       | SW        | 32-bit   | -
// 3'b100 | LBU      | -         | 8-bit    | 零扩展
// 3'b101 | LHU      | -         | 16-bit   | 零扩展
// =============================================================

// =============================================================
// 小端序 (Little-Endian) 存储格式说明
// =============================================================
// RISC-V 采用小端序: 低地址存放低字节
//
// 例: 存储 32'hDEADBEEF 到地址 0x00
//     地址    内容
//     0x00    0xEF  (最低字节, din[7:0])
//     0x01    0xBE  (din[15:8])
//     0x02    0xAD  (din[23:16])
//     0x03    0xDE  (最高字节, din[31:24])
//
// 读取时按相同顺序拼接:
//     dout = {mem[addr+3], mem[addr+2], mem[addr+1], mem[addr]}
//          = {0xDE, 0xAD, 0xBE, 0xEF}
//          = 32'hDEADBEEF
// =============================================================
//
// 初学者提示:
// - {{24{mem[addr][7]}}, mem[addr]}: 把最高位复制 24 次，实现符号扩展
// - 本模块没有做"地址对齐检查"，默认软件会给对齐好的地址
// - LW/SW 地址应 4 字节对齐，LH/SH 地址应 2 字节对齐
// =============================================================

module dm(
    input         clk,        // 时钟
    input         DMWr,       // 写使能
    input  [7:0]  addr,       // 地址 (支持 256 字节)
    input  [31:0] din,        // 写入数据
    input  [2:0]  DMType,     // 访存类型
    output reg [31:0] dout    // 读出数据
);

    // ---------------------------------------------------------
    // 1. 访存类型常量定义 (对应 funct3)
    // ---------------------------------------------------------
    localparam MEM_BYTE   = 3'b000;  // LB/SB: 字节
    localparam MEM_HALF   = 3'b001;  // LH/SH: 半字 (16位)
    localparam MEM_WORD   = 3'b010;  // LW/SW: 字 (32位)
    localparam MEM_BYTE_U = 3'b100;  // LBU: 字节 (零扩展)
    localparam MEM_HALF_U = 3'b101;  // LHU: 半字 (零扩展)

    // ---------------------------------------------------------
    // 2. 存储器定义与初始化
    // ---------------------------------------------------------
    reg [7:0] memory [0:255];  // 256 字节存储空间
    integer idx;

    // 初始化为 0 (用于仿真)
    initial begin
        for (idx = 0; idx < 256; idx = idx + 1)
            memory[idx] = 8'd0;
    end

    // ---------------------------------------------------------
    // 3. 读操作 (组合逻辑)
    // ---------------------------------------------------------
    always @(*) begin
        case(DMType)
            // -------------------------------------------------
            // LB: 读 1 字节，符号扩展到 32 位
            // -------------------------------------------------
            // 将字节的最高位 (bit7) 复制 24 次作为高位
            // 例: 0xFF -> 0xFFFFFFFF (-1)
            //     0x7F -> 0x0000007F (+127)
            MEM_BYTE:
                dout = {{24{memory[addr][7]}}, memory[addr]};

            // -------------------------------------------------
            // LH: 读 2 字节 (半字)，符号扩展到 32 位
            // -------------------------------------------------
            // 小端序: 低地址是低字节
            // 符号位是高字节的 bit7
            MEM_HALF:
                dout = {{16{memory[addr+1][7]}}, memory[addr+1], memory[addr]};

            // -------------------------------------------------
            // LW: 读 4 字节 (字)
            // -------------------------------------------------
            // 小端序拼接: {最高字节, ..., 最低字节}
            MEM_WORD:
                dout = {memory[addr+3], memory[addr+2], memory[addr+1], memory[addr]};

            // -------------------------------------------------
            // LBU: 读 1 字节，零扩展到 32 位
            // -------------------------------------------------
            // 高 24 位补 0
            // 例: 0xFF -> 0x000000FF (+255)
            MEM_BYTE_U:
                dout = {24'b0, memory[addr]};

            // -------------------------------------------------
            // LHU: 读 2 字节 (半字)，零扩展到 32 位
            // -------------------------------------------------
            // 高 16 位补 0
            MEM_HALF_U:
                dout = {16'b0, memory[addr+1], memory[addr]};

            default:
                dout = 32'd0;
        endcase
    end

    // ---------------------------------------------------------
    // 4. 写操作 (时序逻辑)
    // ---------------------------------------------------------
    always @(posedge clk) begin
        if (DMWr) begin
            case(DMType)
                // ---------------------------------------------
                // SB: 写 1 字节
                // ---------------------------------------------
                // 只写入 din 的最低 8 位
                MEM_BYTE:
                    memory[addr] <= din[7:0];

                // ---------------------------------------------
                // SH: 写 2 字节 (半字)
                // ---------------------------------------------
                // 小端序: 低地址存低字节
                MEM_HALF: begin
                    memory[addr]   <= din[7:0];    // 低字节
                    memory[addr+1] <= din[15:8];   // 高字节
                end

                // ---------------------------------------------
                // SW: 写 4 字节 (字)
                // ---------------------------------------------
                // 小端序: 低地址存低字节
                MEM_WORD: begin
                    memory[addr]   <= din[7:0];    // 最低字节
                    memory[addr+1] <= din[15:8];
                    memory[addr+2] <= din[23:16];
                    memory[addr+3] <= din[31:24];  // 最高字节
                end

                // SBU/SHU 不存在，不需要处理
                default: ;
            endcase
        end
    end

endmodule
